module tea

fn test_simple_tea() {
	// part 1
	key := [u8(0x00), 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00,
		0x00, 0x00]
	plain := [u8(0x00), 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00]
	enc := [u8(0x41), 0xea, 0x3a, 0x0a, 0x94, 0xba, 0xa9, 0x40]
	rounds := num_rounds

	mut c := new_cipher_with_rounds(key, rounds) or { panic(err) }
	mut ciphertext := []u8{len: plain.len}
	c.encrypt(mut ciphertext, plain)
	assert enc == ciphertext

	mut plaintext := []u8{len: plain.len}
	c.decrypt(mut plaintext, enc)
	assert plaintext == plain

	// part 2
	key1 := [u8(0xff), 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff]
	plain1 := [u8(0xff), 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff]
	enc1 := [u8(0x31), 0x9b, 0xbe, 0xfb, 0x01, 0x6a, 0xbd, 0xb2]

	mut c1 := new_cipher(key1) or { panic(err) }
	mut ciphertext1 := []u8{len: plain1.len}
	c1.encrypt(mut ciphertext1, plain1)
	assert enc1 == ciphertext1

	mut plaintext1 := []u8{len: plain1.len}
	c1.decrypt(mut plaintext1, enc1)
	assert plaintext1 == plain1

	// part 3
	key2 := [u8(0x00), 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00,
		0x00, 0x00, 0x00]
	plain2 := [u8(0x00), 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00]
	enc2 := [u8(0xed), 0x28, 0x5d, 0xa1, 0x45, 0x5b, 0x33, 0xc1]
	rounds2 := 16

	mut c2 := new_cipher_with_rounds(key2, rounds2) or { panic(err) }
	mut ciphertext2 := []u8{len: plain2.len}
	c2.encrypt(mut ciphertext2, plain2)
	assert enc2 == ciphertext2

	mut plaintext2 := []u8{len: plain2.len}
	c2.decrypt(mut plaintext2, enc2)
	assert plaintext2 == plain2
}

fn test_invalid_key() {
	key := [u8(0x00), 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00,
		0x00] // , 0x00
	c := new_cipher(key) or {
		assert true
		return
	}
	assert false
}
