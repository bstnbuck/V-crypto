module v_crypto
