module salsa20

import encoding.hex

fn test_xsalsa20() {
	rounds := 20

	key0 := hex.decode('0000000000000000000000000000000000000000000000000000000000000000')!
	nonce0 := hex.decode('000000000000000000000000000000000000000000000000')!
	counter0 := u64(277372)
	plain0 := hex.decode('766572792073686f7274206d7367')! // very short msg
	out0 := hex.decode('760649bc45e628ab45ab83f2710f')!

	key1 := hex.decode('0053A6F94C9FF24598EB3E91E4378ADD3083D6297CCF2275C81B6EC11467BA0D')!
	nonce1 := hex.decode('404142434445464748494a4b4c4d4e4f5051525354555658')!
	counter1 := u64(277372)
	plain1 := hex.decode('766572792073686f7274206d7367')! // very short msg
	out1 := hex.decode('d0df8be036e7d95728040244ef2f')!

	key2 := hex.decode('0558ABFE51A4F74A9DF04396E93C8FE23588DB2E81D4277ACD2073C6196CBF12')!
	nonce2 := hex.decode('404142434445464748494a4b4c4d4e4f5051525354555658')!
	plain2 := "Ladies and Gentlemen of the class of '99: If I could offer you only one tip for the future, sunscreen would be it.".bytes()
	out2 := 'b287ce1bea7e43c40f4cf2b87ffb0bf77b1cdf80c6ca09e2ccb12b2c62766ea52d9b8d5c43d4969b55063cee81dcdaf565614e747173f9cbefe8d33e7b6a9a0dc419502788739c40841e6f0bbf533630b8f829d65748bfab487fcb6da50d881b85407ec3694e45be74ac4fb4c1dd654c5b3a'

	key3 := hex.decode('0A5DB00356A9FC4FA2F5489BEE4194E73A8DE03386D92C7FD22578CB1E71C417')!
	nonce3 := hex.decode('c047548266b7c370d33566a2425cbf30d82d1eaf5294109e')!
	counter3 := u64(1)
	plain3 := hex.decode('5468652064686f6c65202870726f6e6f756e6365642022646f6c65222920697320616c736f206b6e6f776e2061732074686520417369617469632077696c6420646f672c2072656420646f672c20616e642077686973746c696e6720646f672e2049742069732061626f7574207468652073697a65206f662061204765726d616e20736865706865726420627574206c6f6f6b73206d6f7265206c696b652061206c6f6e672d6c656767656420666f782e205468697320686967686c7920656c757369766520616e6420736b696c6c6564206a756d70657220697320636c6173736966696564207769746820776f6c7665732c20636f796f7465732c206a61636b616c732c20616e6420666f78657320696e20746865207461786f6e6f6d69632066616d696c792043616e696461652e')!
	out3 := hex.decode('09026430e4e95ef79103694704783beafe2585a3e9fe91fec5339327aa924a1a76334394e8185dbf3a8e7407a483132194aeced84ddbc5b71659fdb044b82d44f7e59004720206c808c7276e6645cc2bcfe17d25d12e260e88d8d285a2e44cf4b2c1009a0c8083640292fb31f706f604b32c00e3335af52121dbd8200375792925da0f7462425df1ff9e26179a25540313aa41e018d18803055d1dd57c0cd9309e0932ae3317d3836cf1460b045f3565569608716629bef54ead4ac83ce636e2fe1f5791d22e0138bd46e1e7579e02afdf262012373ccdb74c1f996185ab7777e4bc1a47f408651f842ebacfe015f6438ade9647cc8ad95e9d6edbf73e0e590e5683bcf1155e63c7ec11e2c394749dc2985738c1b62cb43b2ac8bc1d387fa929b3c8f6688de132ec2d247d153bf8c7e5')!

	key4 := hex.decode('0F62B5085BAE0154A7FA4DA0F34699EC3F92E5388BDE3184D72A7DD02376C91C')!
	nonce4 := hex.decode('404142434445464748494a4b4c4d4e4f5051525354555658')!
	counter4 := u64(4)
	rounds4 := 8
	plain4 := hex.decode('10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001')!
	out4 := hex.decode('e543b0dab98f742edc8d43f829e28d5446bba338d64f9d9975ab9d6e1dc73b1649d119f266fea62a76561d466348021aac156c63a9a1ee13620179aea7a8deae93b4c2de1c5c32e4b2e5167aceef40220197dfc38027cb91dea38d')!

	// test0: check zeroed key + nonce and set_counter
	//
	mut c0 := new_cipher(key0, nonce0)!
	c0.set_counter(counter0)
	mut enc0 := []u8{len: plain0.len}
	c0.xor_key_stream(mut enc0, plain0)
	assert enc0 == out0

	mut dec0 := []u8{len: plain0.len}
	c0.rekey(key0, nonce0, counter0, rounds)!
	c0.xor_key_stream(mut dec0, enc0)
	assert dec0 == plain0

	// test1: check manual encryption/decryption
	//
	mut c1 := new_cipher(key1, nonce1)!
	mut enc1 := []u8{len: plain1.len}
	c1.xor_key_stream(mut enc1, plain1)
	assert enc1 == out1

	mut dec1 := []u8{len: plain1.len}
	c1.rekey(key1, nonce1, 0, rounds)!
	c1.xor_key_stream(mut dec1, enc1)
	assert dec1 == plain1

	// test2: check encryption/decryption function
	//
	enc2 := encrypt(key2, nonce2, plain2)!
	assert enc2.hex() == out2
	dec2 := decrypt(key2, nonce2, enc2)!
	assert dec2 == plain2

	// test3: check encryption/decryption with different counter, rekeying
	//
	mut c3 := new_cipher(key1, nonce1)!
	c3.set_counter(counter1)
	c3.rekey(key3, nonce3, counter3, rounds)!
	mut enc3 := []u8{len: plain3.len}
	c3.xor_key_stream(mut enc3, plain3)
	assert enc3 == out3

	mut dec3 := []u8{len: plain3.len}
	c3.rekey(key3, nonce3, counter3, rounds)!
	c3.xor_key_stream(mut dec3, enc3)
	assert dec3 == plain3

	// test4: check encryption/decryption with different counter and rounds, rekeying
	//
	mut c4 := new_cipher(key4, nonce4)!
	c4.set_counter(counter4)
	c4.rekey(key4, nonce4, counter4, rounds4)!
	mut enc4 := []u8{len: plain4.len}
	c4.xor_key_stream(mut enc4, plain4)
	assert enc4 == out4

	mut dec4 := []u8{len: plain4.len}
	c4.rekey(key4, nonce4, counter4, rounds4)!
	c4.xor_key_stream(mut dec4, enc4)
	assert dec4 == plain4

	key5 := hex.decode('0F62B5085BAE0154A7FA4DA0F34699EC3F92E5388BDE3184D72A7DD02376C91C')!
	nonce5 := hex.decode('404142434445464748494a4b4c4d4e4f5051525354555658')!
	counter5 := u64(18446744073709551014)
	rounds5 := 12
	plain5 := hex.decode('5468652064686f6c65202870726f6e6f756e6365642022646f6c65222920697320616c736f206b6e6f776e2061732074686520417369617469632077696c6420646f672c2072656420646f672c20616e642077686973746c696e6720646f672e2049742069732061626f7574207468652073697a65206f662061204765726d616e20736865706865726420627574206c6f6f6b73206d6f7265206c696b652061206c6f6e672d6c656767656420666f782e205468697320686967686c7920656c757369766520616e6420736b696c6c6564206a756d70657220697320636c6173736966696564207769746820776f6c7665732c20636f796f7465732c206a61636b616c732c20616e6420666f78657320696e20746865207461786f6e6f6d69632066616d696c792043616e696461652e5468652064686f6c65202870726f6e6f756e6365642022646f6c65222920697320616c736f206b6e6f776e2061732074686520417369617469632077696c6420646f672c2072656420646f672c20616e642077686973746c696e6720646f672e2049742069732061626f7574207468652073697a65206f662061204765726d616e20736865706865726420627574206c6f6f6b73206d6f7265206c696b652061206c6f6e672d6c656767656420666f782e205468697320686967686c7920656c757369766520616e6420736b696c6c6564206a756d70657220697320636c6173736966696564207769746820776f6c7665732c20636f796f7465732c206a61636b616c732c20616e6420666f78657320696e20746865207461786f6e6f6d69632066616d696c792043616e696461652e5468652064686f6c65202870726f6e6f756e6365642022646f6c65222920697320616c736f206b6e6f776e2061732074686520417369617469632077696c6420646f672c2072656420646f672c20616e642077686973746c696e6720646f672e2049742069732061626f7574207468652073697a65206f662061204765726d616e20736865706865726420627574206c6f6f6b73206d6f7265206c696b652061206c6f6e672d6c656767656420666f782e205468697320686967686c7920656c757369766520616e6420736b696c6c6564206a756d70657220697320636c6173736966696564207769746820776f6c7665732c20636f796f7465732c206a61636b616c732c20616e6420666f78657320696e20746865207461786f6e6f6d69632066616d696c792043616e696461652e5468652064686f6c65202870726f6e6f756e6365642022646f6c65222920697320616c736f206b6e6f776e2061732074686520417369617469632077696c6420646f672c2072656420646f672c20616e642077686973746c696e6720646f672e2049742069732061626f7574207468652073697a65206f662061204765726d616e20736865706865726420627574206c6f6f6b73206d6f7265206c696b652061206c6f6e672d6c656767656420666f782e205468697320686967686c7920656c757369766520616e6420736b696c6c6564206a756d70657220697320636c6173736966696564207769746820776f6c7665732c20636f796f7465732c206a61636b616c732c20616e6420666f78657320696e20746865207461786f6e6f6d69632066616d696c792043616e696461652e5468652064686f6c65202870726f6e6f756e6365642022646f6c65222920697320616c736f206b6e6f776e2061732074686520417369617469632077696c6420646f672c2072656420646f672c20616e642077686973746c696e6720646f672e2049742069732061626f7574207468652073697a65206f662061204765726d616e20736865706865726420627574206c6f6f6b73206d6f7265206c696b652061206c6f6e672d6c656767656420666f782e205468697320686967686c7920656c757369766520616e6420736b696c6c6564206a756d70657220697320636c6173736966696564207769746820776f6c7665732c20636f796f7465732c206a61636b616c732c20616e6420666f78657320696e20746865207461786f6e6f6d69632066616d696c792043616e696461652e5468652064686f6c65202870726f6e6f756e6365642022646f6c65222920697320616c736f206b6e6f776e2061732074686520417369617469632077696c6420646f672c2072656420646f672c20616e642077686973746c696e6720646f672e2049742069732061626f7574207468652073697a65206f662061204765726d616e20736865706865726420627574206c6f6f6b73206d6f7265206c696b652061206c6f6e672d6c656767656420666f782e205468697320686967686c7920656c757369766520616e6420736b696c6c6564206a756d70657220697320636c6173736966696564207769746820776f6c7665732c20636f796f7465732c206a61636b616c732c20616e6420666f78657320696e20746865207461786f6e6f6d69632066616d696c792043616e696461652e5468652064686f6c65202870726f6e6f756e6365642022646f6c65222920697320616c736f206b6e6f776e2061732074686520417369617469632077696c6420646f672c2072656420646f672c20616e642077686973746c696e6720646f672e2049742069732061626f7574207468652073697a65206f662061204765726d616e20736865706865726420627574206c6f6f6b73206d6f7265206c696b652061206c6f6e672d6c656767656420666f782e205468697320686967686c7920656c757369766520616e6420736b696c6c6564206a756d70657220697320636c6173736966696564207769746820776f6c7665732c20636f796f7465732c206a61636b616c732c20616e6420666f78657320696e20746865207461786f6e6f6d69632066616d696c792043616e696461652e5468652064686f6c65202870726f6e6f756e6365642022646f6c65222920697320616c736f206b6e6f776e2061732074686520417369617469632077696c6420646f672c2072656420646f672c20616e642077686973746c696e6720646f672e2049742069732061626f7574207468652073697a65206f662061204765726d616e20736865706865726420627574206c6f6f6b73206d6f7265206c696b652061206c6f6e672d6c656767656420666f782e205468697320686967686c7920656c757369766520616e6420736b696c6c6564206a756d70657220697320636c6173736966696564207769746820776f6c7665732c20636f796f7465732c206a61636b616c732c20616e6420666f78657320696e20746865207461786f6e6f6d69632066616d696c792043616e696461652e')!
	out5 := hex.decode('d388dbb472faea6163e45792257d3cbbe418e49f60af6c63347623e484b9d380b7589208708d9e781d00d3d7ac2d2f87cdfd83682dea8607f2c5e775aa51945d542aca9cc270a2f054686f3db4a5c485ec1567b2d2d58b9789a30087a34f2782b3c9f76c763c4c237966761a9594eba2c3861ddceaea69a3e9cbe9ea4bcfe047fe35d38b920386732db081f150456dfd2c1762a5a503083c258ceba85073c99775935de9c0e8bace385c75b62cc62d30a511b5a1b39c00f5ebd335b6f03262b42faac4b88acc67ba0c0f2bdde78340e2166eb89cea0e526f6a0eef7b556ad2ee25c2929ced5d4e079bd2e5d241bce2d24e218359a8099d6b8eb8202c4bd3086b9d611d8a42dfe676186a5ee489abdf9ae89c84fdd9c5ca27e719d79a4436c86c926d5f79ade5d3d57a1491bb8740e19cf532591dc4a26993dad28c7e20ca6ff12a0828c36edc28a6d657212f6a46997294a1d1200edf7c27411b444a3cbb1acd963574a614e6b24cadee175369663c1e77aee2ec6baeb54d7cc7668eabe5ca66a43c085a5687663ec2cbef6283b402d0f458b849ebbb32f89eb49835d9e9eb7a9c5b8837de9b3585f4b77f1d9c555576e32f755cfee600eb6fa3568d7b9993c3af159c2ce4eaabc95e3be1d2ba6aba5c7159a57de17236129fa506b33a243e0d7b253b1619d17dbe8ae63d9e2e321a345ae3bb9185b8e0f9294e1ab5c11e63aafd5834e4196c173cbe9bd54bbacbf6a48bfd669a575c26cd1d15961d108759375569496a21a34e0b1e575fd1e5f29e6bfe8800d1ccf5015d39c797705cea573d97a4515a7040c857656a896ab9923a411bfda4c298d0f88024fabd17825459c29877e042ce775ebb0ad3b038b41414b8ca631f042ee1b3821b5a11cc504e3107e42e74fb97c3394414352065121d6a4cd7221c1a037d860368cc9f16365b38d26d9ed97297fa9314725ee6780ab73f6096ac8c324ad8b8054484817613acda7a6eff5303b570b3ca6ca47e6a7332a20b1442c96b9b7f8e5778965505caae20205f056cd1058f6d447cba4105fc1c7cb4d9cc454600cf00f3828139a9972117dd890ef07dbde7c6bb3264771f456583ab26551c1fd2e177c83d8b87e5468faa35a8551883ecfe6cb655db890f6147e36ef12327eed8ab69727fe8d7824279d4a3e4ea521d68d6a318390c1037644784175edb65c8b9e5e82818b8aced0922ed6bb4ac5a9425458d07348f9aa92af78cdb88051a9f04f1437111f76153cfd3d61bb1b02fcee05f7ef422ac899d8173eb8a122e16d4d723069ebd57e9a1b21b699163783057905973de88a374924d6129b6d6958c6a7d6404007ad49ccf6108c0f9899febeefca32393951a5b49e8ebe43ada86999c1bfb71e38cd1a1f1fae991ecf5eb11a66a5ca8c52e25004c72c847a6f395ef9b6a93bfc51af7035a18f2889ef3eb06596d62f15bd43cb1a024802a71615c46274507d587dead50b0f62794df80cdf68fc9208ba730d508f8f1ef114ef8098d3c7adca8de3adcfcd9c37e96d22d1e9402265d806df1ad285f447435adeae46124bb79c760c90a9e6a555ba0acec8f025919d4d79ba40dcfe7acebf7fb3859c97ea308cafc35792d98738a80ebc78387be9b7604fb53cbe29e48aa5f454a864a48ccefea734deebc089dca2ec8a4cb78fd6d32dbe9cfe097590efb198970919825d0ff016f000a2a45f6365c2f6375a203a95b744ff129c5798247c11aea15a4770e94cd2751787a3751827578e0831013a08e6e4efa9dc3191a4dbe3fd324bc5040e7de896004e3ddb9965eb46832a53a4ce51902263aa1b05a0510466fda753ec5aab1af150243176083cf640b2c385e20a0620f5b13360ecd71e4260014811176b725fbbafe829e420b528c49d978b1c29b05e8c60e173aaee871e57815c0abdaf1bc919f3082d6c6d8a5f9ac029226e894bd9026c0dccfd964b9abe954de1e819c798ef1c5ad32226596e300d3e033161857433d7877a9168aad16812f8fe7aa23cb088ee067f7e95e3c29c23b89a2fc64118738c66e3403667e8fae401bc76aea24870cf09e7696427416615bc5d8dabb5e4d414d65c2e85b198eeafb96b33c8b45750715542b3f985ed00a0b164befca12a50c23b29ec01e576eca5369d5076382a45b6a2dc7f9aad50054e58c2083ecf69d662f0a014c9e615d14b913a6d8913ab50a7e299c92b1f7b5f5c7d7128b77c33b15e9cafe2730da39941fbd58b3a0741752f210b8a49c9fa5ddbc26810e43b4f12fe4afa460d1cd5ab77ec7fa1e8b02cf4e274088903396c3e117174802a5838c8c3e2c7cadf01a1f06b43d7aaf36bc40c3e66d8cd7d899d1379d3a45b41a8d48efdf7062eac4beeabb7a76e5a967fe8884acd67ec9b115db3f43b3e615988cefd42fcda9c6b3211ef3013f5dd4370db52e74ed64f810a7192a8776dbc68ae446d8abcd89c9b2892b81f1dee34c50286802256d34121c3e4df2b2fb210e04b2205aba022e3c23d7466498e73c56680ca88c9c9e8edefa5bf9774c00c624fbad7f230991b2b594d94faf71c57effccac57fc845a65114bb37eaa2c9d2862d365f8201eb6c52acd98ca1051183e463f0717047379d4f3182be975c0712e59b1ec686b95703844b0ddceec583b563fb14108443e03933ab2fbe47c0b3c08c58b0b558d23581f2a353388042326da14db3b4de244649d308bc898287812887722c36ffc506e7e6c9c05af76934436681a6dd19eba4df5411e5ce9129a37eed0074d15916a16e25130bb552f710cb2ad2724502e6adff8c52e3668e882dda0fe7f5722f7b904bd15cb3da80e3ddb720b5413a8251c752e212eec98d2a06373c483d425d49f4319a77f58ead3af530cee9267ecb3cd49e6ae0b2248576d69382c9c80dea0031e6185ece3b2e7719cd5c48756ff600f7f0d3769a9302164571203bee9b3ca3a39ebf0ad2bff92e49614f8b8013649da13245f86dae96fa031fd4bad1b23af789650dd9780e2813975f9723dcc5c9431425c8090b11776c2ce6d63b79a8172588ec1f76c19e8b9b400ada9f59bc0349d0321b838e813b37e306d6ced5e9210de4a64001b4b64fcefeeaf22431b51a78b3977b6b7af45f916c7796a0184500bc504ec379d442db3d99b09dc693fbbea4c2b4646cf81b3d7d10ef22f3ba72fa61d97bbc2b41c509d01bdaf771df109d3fe8d62fe438c82e6f8d0f5fb8a238e56982082b4c89196933c2fc02b9541574dba8a5ed568a61dd0200fd6df4cdb1ac22e2c07eb5cc94dec0a3aa5427483e6f1005b4db4f49eabf5d730db212a18b17d2b957a15819f502cae22b3f3d6c8fb0e91e36e67b47d9f31a45bd28926efa566fcabc9fd680cd14c9eb5f6b5fc864f9774359d6702822f43d947573724fcfd605b876da5aa82c843c7fa04df45f046cfd62727c70d7dee')!

	// test5: check encryption/decryption with with high counter value and 12 rounds with big input
	// out5 is not fully approved for correctness!
	//
	mut c5 := new_cipher(key5, nonce5)!
	c5.set_counter(counter5)
	c5.rekey(key5, nonce5, counter5, rounds5)!
	mut enc5 := []u8{len: plain5.len}
	c5.xor_key_stream(mut enc5, plain5)
	assert enc5.hex() == out5.hex()

	mut dec5 := []u8{len: plain5.len}
	c5.rekey(key5, nonce5, counter5, rounds5)!
	c5.xor_key_stream(mut dec5, enc5)
	assert dec5 == plain5
}
